VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO GF180_RAM_512x32
  CLASS BLOCK ;
  FOREIGN GF180_RAM_512x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.000 BY 1.000 ;
END GF180_RAM_512x32
END LIBRARY

